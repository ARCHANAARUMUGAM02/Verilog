`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.07.2025 11:15:58
// Design Name: 
// Module Name: binarytogrey_df
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module binarytogrey_df(input[3:0]b,output [3:0]g);
assign g[0]=b[0]^b[1];
assign g[1]=b[1]^b[2];
assign g[2]=b[2]^b[3];
assign g[3]=b[3];
endmodule
